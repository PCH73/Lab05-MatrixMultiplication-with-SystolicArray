//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//      (C) Copyright NCTU OASIS Lab      
//            All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2022 ICLAB fall Course
//   Lab05			: SRAM, Matrix Multiplication with Systolic Array
//   Author         : Jia Fu-Tsao (jiafutsao.ee10g@nctu.edu.tw)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : TESTBED.v
//   Module Name : TESTBED
//   Release version : v1.0
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################
`ifdef RTL
	`timescale 1ns/10ps
	`include "MMSA.v"
	`define CYCLE_TIME 20.0
`endif
`ifdef GATE
	`timescale 1ns/10ps
	`include "MMSA_SYN.v"
	`define CYCLE_TIME 20.0
`endif

module PATTERN(
// output signals
    clk,
    rst_n,
    in_valid,
	in_valid2,
    matrix,
    matrix_size,
    i_mat_idx, 
    w_mat_idx,
// input signals
    out_valid,
    out_value
);
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
dSbxA0mwQOrahGKVqMhdn1cm+cBH1PBhKnYd6XKlrBKPkAECBnf+XfO07HQSyjUR
XjOwEVtZ3rLDAJ9HGB+HgBDxyQEJUc67DVxWb3w3hBkWg35iv3QzEnHK2k66lfBA
FJK/A/6ZE3J2YxFRXZcNh5n6alNn7h/ZSDRf8lJVOSMrcMqSYqfaEA==
//pragma protect end_key_block
//pragma protect digest_block
04fRGGtzYzxWSd00dsOrCsOkbkg=
//pragma protect end_digest_block
//pragma protect data_block
f4hfRKdnaqpxNAw7FWDLZozu95q0Moo29y6lveipW9CctD9g4yygWZhJEPYTJCLd
rQDfDBpBXyCdfBrNQSEZ2rZcQWPS8QtFNwS2DPFn1KmCoSWc77Z8Giq0FBitZw4K
WJnrxbXq9vCWeSTAKHlA2qhAMjbltLtCr48zBI88EfZnrObOzDXYUJVGTq9fmilS
jOUodvEPa2r6Uh927VQ+9kFkb0L1FUNyUpkF3B23x0iqROhEaYsk1A0N5W6b8j+T
9py1Q/+MNGTJN5PPk7zB1oluHE3F9ecXe15ifFUFZklUdaPQfXBvPJ+krOjAxFoQ
uM3Vh0qIRKetLqnpMwOB4Yo/z24Son49TL7qwlVMoit3Hb4gFDdw3Lth4/vuzPa9
PfSTjX6NcL8Fd43amQWenGrAZQxDQD9rpTL9YL/pjQZ843csAOla6WqA3bnSoaLi
2SGSGX3XTYGymnMQGTbjfH8Xe9cwYpmQtKehHBU0xerU4Y1pCi5uvuyYdEwkxFFl
rXCqJF0W6Z+ZI0/LylQs7VMD8zfdf/sdCvY1GsRq9nj3hFOtbPTR+kvaEaprTTtc
eV8tSGE7r0na9DHArXOliwsYDfsG4fJ25Ft17zZxQu0+tn8PXzILn36XZu/IvhMY
A/cCRIj6r6qd6KSitzln1EX8KLGIiEeW1Sv7HBG97eOCAVRaK2HqStP+oPjxDvLF
cavKzZyuMeIGZfBPmM5lYlskK/jH5uhkqbbtU/NqIUJkiYl2tANUOPT7WLfDCft/
j01BTCUthkfezyQ0F8UOkmWu42WpsSrBk06x5vWrU/COEQTJpTl/jlF7ApKI8zf4
LSVRFjFLZtHUpplJjpZnoYryXh+a3mhssC0/rmtEs7P8CMFFXvBAQMajp5dlLmEt
sFsTPHffxnB9gVZxXTNqtkLnJOqG9deCP6GntAlOHQ7X9qnSxJxUY8hGIR08MykZ
daIdiltVxUrufRzRDUz5qDCV36wBJxKTChwDOSBcqm0YX8ndVVwv8u0ZyvmXVysX
pziERDWvKXT0lgN3DW1RqA6jo/7BHix1mPuhLatvWS5mZ56H1nQj52jGr+9NLiHR
/uQqjChsGm/934AD8iwcj7VhXT3twpCg0BAx/LONw16Ug0YTiBO55hcg5JICDPEs
MAUI7trIn3HoIP8zYbkBpPsnl6vnijAAUxPkf8DvEOVsk4JwfgXhDfhwqnv7iChR
MInGhuEjN7XboaVNjipO+pHg1QHIeMNRcvTpJbG26VfvUz85eElIxJtsSdxn88Aj
Ou38H5GshBslEb8PjSDz8KZ/oZv+HFUmgJXgdzS1h/xNJ3d98cx1ytSkW3RNDZCm
f50nxPP8JT9LIQvhrUT46aSO7+YmrN2EVcnJFe5UvQVkBtKqvYED3skVo/9OFWqz
YYtwqlm4mFhEteQ2/pP9JxDsh2LCg9ptNGX2EW3cM06Q23kt8Eo/4jghLvyille6
el7amYeqBCfpd0nu2Y6lYP6LWXqJ9zneUzf3WXhFE2642kbIL/tYBQNVFUr5jblh
CfUV4dSXunVhcKeUFInBDdj70RWuLgWFO1t6CDovZgcLpcFHRPqPzuaRcdRSH2cf
u4tlFGfyBp03rhgJvHyN9PdmCofVpwO/IuOP7cvTrQhDdhVAwqQpwP3oW8rG7VGY
/sShUPYi0fEQWezspxiaVkdHG8yoPSMilOgq34G6FJltCnhs+bkE1/l5RYfNL/Ul
TGkUIodDVHWzPDlDUcK9VWDKnzXUaRE5VwCUOnHknOwEwIMXdlHG78x/Sx9AhLGX
U9x5lUvm6U4qouJcCsbKcFfAuDmKg+YbM/ZtjfFAZFU6QtOyMwRS/LSKURzH6eAG
2PTUYDaMSviFxRHjjApQNJavzxySSFPP3F/yf+b8QHeASrQbcm1nVgLZ3U/fJ91L
GDz5QP3tBF9ifY/NDFLxrwj6h5lP/TnqZrfySdmIGwbf4k1acOUuAtJXtXhXTc89
rZtWnA6Pi5X8wf48uSH4NYhidoicWDEx8Ilh9WGxnaWdiOW2ekqjYzox1odAsMir
gHx1jNwDBQFygrx27y3zZhHBGbOCgwdBuF9xtiXpPlgeEHXf5rJt9JeV/pV7xccY
O7MF3gjhfxn9kH/+le5/WCzhQsV3eKG1bfpkJ7YJchMo12bkKnEp4NO+49AKAwth
RVEoqnyWcNlISHGw143QP2nWWKGvTf9CikYItl9hIuy6YElbRvpZMgr2X76iEiHd
NuqTH6RSCghr53YR04eQYJGoRqel+HriSwXsF5d/dt9AIKWaJ6wh3480qZmDcuDx
ab8/4K8aayVSteMWjzgnYm4na0hrLKHi20gpkKSQj0LXybrYNWr67UKfn81tf/Py
Mx9qihIjpF/bzspLQdjDMbTl4LDOq7mG2DK4n1/bRmGyYW0RedBjOXMtcBv+D3g7
l9iUfJC/R3u2vy9oq4SyvIguWFSyFCLKQoLyVBhi+Hfuo3DCoUesmdH7dueI1brG
gDXVN/o1OwnxMBJWEhhCZqr8wgM+Y2I4JtUbAh2TVUw1ITvSwtW1GC9hTSH3BdIC
TtnQ+VOzgGYsRxmNJt5pTqb+ssyMslwlvbyLglAH9WlZcFN6dhYUv+QBg4W97wPR
nVRWuuv1N4CEwjjw8Tc5gSV05FAjr2rXk+wALo3a0I5ELaGiVx1kh1Z9+Eysh5Nv
Rh0CyZfJZRtgxuTl/r+pUBF+7sJVMW/g+JZA67xZIXcZHvdk2mQr/0L+dQFOfHf7
y7uKVaJ1NlZf+d2eV3qrl8DLChUXybJnFsr16MYPYOJdqUxPATN6lt0u5uEN7Uwl
VDqqP18N4vw5YUgab1pN+rLJBOlIaLfFZqx9dyjpuL65emNz/gprwikAuaqQlYiX
Bs3DLKlgfldF7xcobNzcNw1qvuSe8aNYF4Ycu+O7eTbc8kfjmspRp0ZE7LhR0y87
qzYG17ky+eVedN+mQPrMbV9nnQ2i+pllgNU+NAmcePIBe6p0pxLx1/KDzkTyD4Yp
mMhxszTatDW06qc31si6RhF34m66VG4rvs/mIFZ0Uz6gPgcIl8q2FYkVNh5nH+l8
OAe60Prv9k8zihzaPLHrgtlCf2U3FWQGS9jsJmFg37AhpCxQE9+uyO7Xa2lu7fv6
alhe4j/G8WdaJ8JkCiodws93BN1WN0NzULcu1oDLuqHDBSobYC9+3WzGPGWrxrqQ
fLGWZh/oWk/rDSCxZjDjjcdtyCuFc5WhKKzApg7tQDYkYlcj8XDaw4sTmCasHhKk
nxTm32nGRziamRgq4ZgWsCQMAEBvY1iUTz/jj1YFOAsT2RY1h64CNI4Rv142G7xn
1jbpuFOGJDAqDDKV6loT6dykbBXQx4HIx4+XHYcKMCn4pItoqkjnTG8fupk7AmwU
HnY9lwv5hzuHZVC/eD2lSs94DmYHm6jKtVYjm58lGPSG0lIAsWUwA/isYtS5iRt/
r8ozrhNV38wHv6XTKTvJUi+uucneKWQp0IrpMbT9y7341D1lrmhZ57xfpS1XmbEu
YOWjnrzDjtFlC5tc3GBLkIe1ZgjugQs6rmKbDacZ6c7AAarPllowhae6+BdJqXAJ
5UWu2xqgS2ghlcw1FH1c1/mbscfPl1jISOazwcS3favP/lwue5+ZCr/btCGJaiIT
yWEgPrNbwsuiVit1HGjahiCXjI7iVCGDBLpgddJuds0AgCqqyRg4pRBoPjcZr163
4cR6S/h0X+7dpb+2PTKePuvM9SRN5FJQ48fpsFNU9QcvYI1TvMVg57bugEQ7AXdP
kRuD+A8bA9QUHIpsvO/UtszWx3Yvb6MV4l8iE2SJQLy2TqES7Z+8oB2vUvEw+37t
1Z/UfMK/ND1v5DgelDK/yBnupv4hwFkBk1tz2rh4QRi14J/VMQnmKk2xH0S8SBYX
cQp8acgQSFJfVIBXMj/v9Sv93D+rPlqneL7e5TZmFY8CSM/QAmQXAiZdLJiIxfJ8
BGtg6aIPKBf0F+4tNQbnvdy2X833vPEJJAD/kpAwts112nDx1wERpjQvFsqIIvXF
uvcWQs6z03SgICKJYZcP1d/0ZvZLfioGEWfSco76C5F9Bz6jxRmeP4Fk91yEGeMS
6ryOx0yE9VD+l941uG57ngY1slR1TD5E7BwxluzToycYOwYjIpQTkK1ow0i6Wnno
2LkK3P6bRfEZDclBWicXmha3G8pfPLK6tC+0RNMd7Wf0XN5tnkO5R0EsSO+EyRTn
nLOAm1iaRFNcpmFtb0mLv46OmYEhSS2ZaUgRmwtFglw6ufPZC9RLWI1ucV4HcTW6
ehBadxI51TDPpE4EFimqz5P5R+LKc9jEX/WWBUh+LEic3mWSdfL4YIunvZq43gPO
KUNvbZ2wbguLWkNYHYhiamrHD996oM+sGUVHctOExi6i5iedGaUT9HF8kdpSH4XW
LZl8acc8hxUvYuK1o+rDE4P2kvFjfXt6g/m3uNwbFtJ28StEKV2x89aTS9TzU6qC
07QCyPv9QQgmN+uewCEtAJip5i9Zenb5pJD6cwD5LVRJGrtnoguB3ZSZ/pQvCufU
BwI1uJQjgW1YFw5OKkgmbe5DLG/0kKci3qFc3+Km0Hflt0ju/N+W+Ap72ZhETCc7
k9CbBPGdN4Poyh5l7KxdrlvlMAStE6wPDbkDAujWivJRPe1jlUexZZoDdEEYLQdA
kUKF//zngxxPzjPZxIZKKaCw5vjNl/beNpfZr/1dmpNVFyiixS4Z0TKqgWC8WMuf
7I2sSwvO+MwXFKnNYnWfqX6ZwY4zIX/Jz21rQMI3Ay4BXWqAPNOG8i8ZHOsAga+L
Yl21eL2wv8sFGuyJgWWEekmLQMMHqGA7mNAbQIBAP5zhkNVImQekF13601msXo7f
cXqLpK+O9pbZFSPSnS7FcAuM7kLvPRD4VIwIxL7B/Pt5J7gob4VLA668RlVSGCGY
yScaR0ijQ6DrgxrHzDeZxZxDZn9XNFuUSjHV3nzZfqHsaKNfmLOPdfhDT4bs9ja9
v+hxw9+9ay6/gBOy+Xrgk0CM0oZPBKUVKn3/g0of6ECcJlPC2MSieRT3TabfJx+A
gh4ne1FCeJc9RqXWC7qtXnpGbxS6DjGmCkK//8fRW1yW90ZmHwlEXyScawAJLnhT
73PEXFxRzrizJezdqhQmiGE32WDtpeQxf1kq7km76iH4lCZZxVDfkhqBnlURMCGn
5AWjpBD87oVNE7OskpV6t978x0MMFYmpJGw6nI58YjtdDCNh8iOsefzmy1U5V6CT
3mUk9KaSOYQILL5FhwJpQ8JzakLYLfAUrBZGXs9tUCPkQvb7HqoFqylwv94lUePd
eLMufrvnKSRmhR6hEyeC9TAUHCmf8YSsUwT1l1AIMHHep7mTvDY5wc4TKpCWXJdm
LaX5hHI4jFyQXgmcfYg2MOlQ7vsvuuUioV6LLiUe38+86fqnf90iwglrTEWET4/m
x+lc3oKX2PNEFC0b60pNiQCC/Y+Gny3wtEq3BpcEKh84MopnEQR49MPVs0ucV2uv
j8bRDOlRjBKSvsh/FwqNqZZTC6KgYGClTLJQTSpeD2hTLsaEDf8hnmVHGugpZPPr
Lr6X5hGAZEphPrf5L2aYrybgdNGGP06Uo4Jp1RAqqBr0BCZJ/EvRLYgVg8AEu+EF
d0e9+xXteBprSCLx66yIBagVlIoOhZfULDVsljAW9Z4YfyXpxhBd4d4cCyHmxQtX
P95RhIjP6Y8eM5JKctdIZfeSJSbslwcBs3ehNBSC2atA+Q8jsyd/QK3JvpS2ZPZr
L8V/iA+CZShrkPElP2uEtBj+qJaVVRperhYsd3aPLMqA4WzhP0D3u5h/JTzMYm11
viLe3UtBC8Ovka89VcTgf7hruU8WpVbPFt/woPQZ/7rrNb0/6dPoZ+k17tMAC4/x
MDOgDlonKV9p9ExB64bRwWoG1EtuEUir8xn5h5nV4G/5/IyHsYO+8qriFY0hY355
5arCMlXB4442ZAEiLswiMFXGu9SbWrkCxtazB5VA44pAI3HmYI9ndUgM6ErS7WrL
F1Nvw/rmU3slbhJyv8uhK0DbD2oNyu/rcgohXTaWUPgMHU4jNyi3hcG8LdnL40Be
mh5TqSkNdn5oqaXWCviQHwr3GigCVZEPBV4VSeCok8AuN5dl+zfyGx5zgS5gBMQB
NxkvlWSGih3gA4Yseo5bxDdYxPwP6Gwy7e9s3Rq1u3ZVkfCi2l44QQauJk3yXaK1
n45iCOqlU+6vDB+AwD12dWJ6A/vMA9u7yC5lSw29hIQlMYKE8r5eNE5YTaRU8kOb
kUsUkSLqXn4HgvboeycSleMN9ZpX/n5ZPtCqEmiUGyufRESafRcP9GxIZkgqP9Cv
IPD3xZx3QyJ2pfXtHwOL2UvUrWnG78aWhsYbGLLNRIHVkLVS2ATVwXRIbSlE+8OT
lA1QarKKc7wLrXHguHMioz2hGEQt7Jz31gTbvGhsT+S5I5t/nFci9/9ze9h5qKfZ
CTt19G6k3Hweh0cCe9IR0Ve6ts7SiD4C0iQC8OylswJJtAnfmjPrNG4BCTFfDb7C
RP+sSKKZE3CNPTJPtfpAsM1qZjLdahWHhu3gTCoIh1BfXsu+xhMifHVwMyc809bq
FhERv/4HDpKu0N4+QdRdD0G/aigQagGATgrchah6QGbrixIQ9LGt2VeKvVexSzjN
wyfYkibIDIY7uk0cR21Rc1T3QWGktBZQ1mPwSxlgHBOafwAztMvwUHnau0LIYQ4P
pC/5F//ks05unkM/zcgDjsyxV7xkU7MS7RDmMUMGeh8pQXGXLqvCsYorxURh2yIk
yxvHo5PPrRw92HFVW6vCfiGCFkl6go6osQVbegvafNbfZ7jaFTvr9hBiQSsY0pfI
GeOaIWBZXo9RwojIohXDWKL6ZzbhMO74BfalPrg0peELUT2wYatof1rL6Jw6o+Gd
KVaXtb04CjlCth3Gk6JdfA57qKl+WhJBL32JrGqr4kaBZ+Onhj9qk7Xo0E58I0cw
rkDuKBTEiyVV4S76dI5LqBlUQVwnwoMhzsD8ncAYJbi6Yc2lPZScsaH3r/f8aTHs
Le6uDmUfG/SXtZqsr6q3T9cyGmepx8jaDTN4MXI7h7i0tjf0SFOL6U0uA9XNlJrG
4Gz8SCCgiP9KkxVmsgWnqMK5HjseC6Ttntf1mP1gtKaOpZx6t0PYwBBIl5LIMW0k
MGPTvVD0f+x2/pB8Nv/6DRHitwHQzu30YltPyEKPhdSQlRpf5SnDRg7j0y6iDrH0
N5sz/6MbHL8BpqmFSHLe+3LbuZBw4i4Bw2IMUeyJfTC5yFLUeDork+wpW/1DMkU6
jhNM4x4taBhtItG9hfPQxTdvMqVQiOOKUsWJvSYOmd24JNnlwr5KtHH1VVXUKlal
Lr89Xu8gGXGOolWeFqfnDIF+JK2kMgVNfQFab76y8FiPjbjsxTts6GqLGhI2eE8N
GofhE+iQX024y/XNPTuzKW2JwOZc39d57JpzKl41b1G8ZohDQ8A4JG40zBqMbscT
KKb1A3piz7attYNw8RlhMPl7Q8AD0pgghSFcd5Bx3BZ8lz8PJ2FjYyn45SSj9Qvo
DoEQPKd6QIRabU+UrxZf3BxO5UA7bumLIk2Vmva1zgKvqB7eNTJzDSnptSLw2dPh
y7yDyU9LrUNh4wFsg+sl8aILRzRceHcOi52+3CZmEBAgb6wAKqQ1v/bAw/Rpj5xp
pmlJSjTMuevCYV3a9dk2yK5d/AMWtF4kT+QwqwXoSGWPaZi2HXntH3O9RLgWZdhX
QdNSLglrMAew0m8pCYYPXEfdlVQUa+94hN5wlPK1zlUZu2lhzS0me/ul2nvfN1En
/LxLxr6egCxCL1rTTmTc1ywceEt13Gx0D+NwNiCIc/IVCMYjLXZ6/0ru1B4YsJWr
01slHQ8zlNMoswS5JA2Qmh9rWapTcTbS+fyz/go7mGOPMr8Ker9s6gJ8lyIliDBc
mVdejTueJ7QcQhsFKnLylbfuwF8omPBop3/Kt7+mU+NvLfNZrpNqO3tSul3Iswc4
juTbUa0f4AaJ5yvTAhWcXX1MqWr7ze2IUPbKeZiPZskH+G1EUWvrcDWxfUEYyOsI
/TvUi4OuTcKn7a8jXyhuO+nVdZ5YQo/oiM+hYXn8I9cn7T9EOS8bJ6IOtm2UgdrF
8FsuueAjs1LGUfS3jGZV2mHnqUA+4vPJbqw/5KsfMbvhQf/J1+BYhh7vd1pzaalP
iCdzBPo8c1hWfS15Ecq0a3hB39fg5rXSRfVWU2udkz5CZf5HNOiIg7J38wUtCFic
LcfilFI5AC0SApAyDrdeMcFmaeVt4Xrl8I4Bh+urwcRatUlD8PVwVNdkBykSJeOp
EBEzU8Qbg924Q+Sncsp43xf9Udr38s2CE/2mCIAHJLLjI+2O5V+wGel/npeBlf5c
aUQhuGNsWEI45NPq7h8I1Fx4hW4G4003O0zxgmoh37+E7lwAckA9qcBAvxab9WZL
9Szm8p+whDpKVoYRid8VRpUsYeBzTiGsumrSwLQMpSdjAgf5MnpPTZJ/jwj6jL5k
TmHQsQbiGs+6WCELJWIF0Q6lp3/5sVwzFhCfhUm2NteX+9HB3WJ5PPHUz5CSaREM
ey9rRJjYxYUvKLe2HdzHNz8tXrLohqlw+eRheDS0rv7gQtJItuvaDwxiDwxye0Lx
Lw+xpAu+q/adiNLoJZk5ZwWCVNsGmwQqb6+TbGrMUvU8xpk6z+gX9xDtFmiNar72
zGC95WH0blXM1GYWzON3kEUVeCPWJ4eplozzTZhlNrjlbKLX3I2Ws/CjuCUATxYT
7qVuajutKCl0mV+K6V7dVkay9Hknrg5gVLr3bPcPWrDM1K3FGDKEsUInCNzEXvOy
dhMZTXycKYJIimi26jBFq8Vv/VXVsOkjR5rmkgBjEg6E2liBHM067/awjGebbcrr
S76e8tkyDJJe4koTd/jLyga0xLSQKJ9jkGjFaOrl66o37J/ylS9eKIQOMVWuZMU1
vp1UfojNpjlASHNLxNquX88wGT+Wtwn0iA+egM89zx54SUyKhFhBoKvqa+AEFHu/
0UZ2EYau2Kagp/97+9u7xN/q86wrwDNt3Nh44EWu/kW/F6N61sI4E5DXlmxjKc8R
ItLnXtXXE4aEOspcRU2Fo4Mqk3/VuiNQsRQYPtimQS3Opid+blrEjH1Tpls3QF6r
5BD53UtFe8FmHs6YbzSFHmhCiz0Spjkp5R+nkXzHnSf1yrz4aBVxGM+AysBtXr9T
euK0YdXnJVPTanW9CuJWzmGKsSbPNg7Heovsdjqu/KUatTbgWdeqhvsqNRUCMPHH
79U7LNsHVXCNh5CIZexdXv14dxXuDkB35JA37zeDxMvz/eM8mRaz16Y5LbaOxeoG
hWW1tUOfDMdScklno5ZGEJ1XRGdiq/EW4KsLJIAcspEXRXDeR2anqVmw/kspkNTm
qkubFyjnP5BLe790UAMCauswlAi1VCSM6kB4ctBa5L9y8RByoN2DzKICMwHTZJV2
YRMRzBktuMoTdhkEv02nA3BQ1GioS/vEvbjfn5BJ/9Yn4fLzLftE85rcIsXCEO5U
EQInqq9LVb4aW4L7FerTDNs/BSLcIn8eHzLY4lDH1J7mUdxvQZAKAoeNA4SsXTnO
RZseLh2rANLZ6TiDOYIjfiIwfMUVeM/8n+cC/0oN+fw/+QcTh8DCUAdVV7lht81K
UsAdQii0lrk5QYMj4rTEaUOH2oJFSl8BqWLbYUbEStB+RXS6G63t2BiMr5WcRBuA
hssAmLzNdzm/OxugDnp6YhoudRoJKSrUU1Z3yawuOSl/pdk7I+ZevLLu8Y+kT7tY
NBpM4jyWhy/O+H/1yekwyAONo7DYO4sDZU2B1z330skrp8W5QsDWTQwK5mIm9JZ1
u70zxGtGM20UQrhKo65dXgB3fPDpl4jCYut3UwrWc+41Y3KIsxU/AeeDHJ9TkSka
O8RysLrSNovK3a4uryuLBdKphXFKt5dAGqDuGsvdfczcrEJJLmfQEw0mucJSO81n
xwz+hdJFoW/YPdCzzvsDIPJMserHGwEAYx4RYF9lxIhdG/U0mR76giVMCYuP4S6O
U2aGR8xLGB6SwD5w2AjxQewQaHTe0/bpYWGKpxLzClDRPLWDnTAd13JEc+r2LahQ
+BwwX8JL2TZ9IqRpg+i9w7UQYcmZTupV2eTZMfxjeCvI8DkFp91QcitCbMRIx1pb
l89XGGzp6jCImhjiPhScivu8q1WXe9qnPdVftiPDoDBPGwTP2LphpG+gfs17O1fu
62QLrYQPrmNHD7RnOv20vA3BtRsSfjH723xNAC8zcFDfXx0bFRj9wb5GAxbW+OK6
RCoKZOAGCW6+76DBkv5TQyvUJUSmYksqDFfJGg92oNVjGV7VN7+Jkh7oblZ/zoPR
HlowaxDS9YeklyUwIJRqBdpj2IEFmTb4tfbrSzyDy/nhJjOzYZZW87fU4G2z+iCi
vCgsmAb+ww/EfIHjnPddf7cbglHjbmwddua5sZndW4YJgMSO2JSIl/3mf7EBBmv/
U1j8kcFAdKSokvl2cHLZb/A59meNnCNsoqwdVqHc+5H9B8+0/5KDZB5jvv5tdC6L
phYX1Q0aXyCkQciN3DHmzu4BXd43O9kKpTXyOnjbu0vZK0DcGCccSuOKhUNKb60h
Kn6gsHbui0imtw3N38SAWOzkUVf7G0V01sFCjsrFGoj8BVhnGo3W4m59wnDrn/54
2+rAtiHzww+zfvfZEp0oDQkW6BZ8w5Yg+c/lhIAOIJM32kEqug2IHyLtkubAH6J2
dea+FJoFwfiU80U51HUJm1lY4Gta5QG7BlUKtYdIFK8obcuT549Ek1ikdH2xp9JJ
BKssunaDUyl392LlOgLfZ4Ef0dB1um4xAk72FAYMBOtSQk2M9998YyBeAH0r9xuw
5y60P6LCZYN0pz3hqVDVUxjr8y1R4on43Cj4oddcYrr1UCLlVN0i1YXPA7U5Whas
o47MrEBnO7svZgwoxyn2YRx/2b3c/J7dTMuFqgAVnYwpvOfILidSTR0QTZdWWIjg
6jwLgTWZKoc9w7guDlh2Fd9Mo4/plK/1w/xanMpZsB9SAYCYjfAop+Puk0sQx7V6
xZCIcLYzoJ8t3kuwN0Atx/JG0m753oqMXCQXdGkFJGFw5KeXiEAUPmLcKzJHSU3q
iBwYOvOy/sbc2pCZz1XAblh6KSh3e0GZz7hyOmmATuF4R/u22x7mINW43+IU3bEE
cG2/nhKe+mWcw1CNumNu8HZ+YzjVx8Lu0V4cqrZJ6con6RDzhkpprLyXbmkE2EKd
htDFofiTDuzdUKGz44DpLfF/Vpz/fG8ciu26JUSjltA31QJN22l0ddaY7qNwPAh9
neOqi2Y8aeVHT9bxrmg9q/6LXvUP9OT1l9UhlmF2wBWkO05e5HYuLGZHR8O9HVRa
dA/THu1a6TdTGA/oWy3h5QXsUDSYMYG1ZScusoMggL+8Z9kDNZhxiP5qTOo7vDhe
jY5lOZ3WL6+bZejQUk/s2SPkEGxSsOCsc+Q/YUPIjA/yr68CVg9OwEeIecpG2fu4
9ztgMWJin6GOjOcMr8cjyTGV7QkifaM7454g3WXAePEnNinmV0QfL1ajMwLlEsj+
1kQKFCArzOF/AsuieOMQJGciRTGF7MiY9a+IkmfvU+tm64rS8vc/EtW+jLmIr28k
Ob73uJwgRjWN5HrcRCeLmvg6vm3ASiZF6/M27877vlCDTub4GO20GTvPWI7wM1qU
EXBeafSx6bDrM8OZoxpJ9de6GlC/rUaaLdhYtMGkmiNgWjqsJdRrWCBvpen+7uA/
5iGRzl4j23PPaE61q4Qc6FtO3YmSKAB9zkPI+kIGEdpIFYs02xLjYTRgl01IenxZ
UwFJmAdGpOhA8zEXbsw8d6UHp+4Mh1oeCD1Uo+DIp7cxzHjZu2F9vMohnPOYhx5i
f3fDswFOWDEa3j23b8+R6/C46PCfJEOzKC6IuH6iJIdBN7P4g7coECXlNTEjrf/U
Z4UxzuxaO4uGpmmFVE7tYa+derlXo6gZ5BriuvwJu3xEgCDDyuanmg0OzLanp1Zm
AXYzVr0EDR5S5WtfyPTOMZ8x4ur/8HS/UZLHG+DFx9CssipgwUh2XZCkdj3JUKGH
2ZH9hdZR8H9AWR1i1tPDez+3drGFgRUWjpu0nf524O2MTpjjeLqfmJdUgmUcvyHP
TEfE41umUAL6mHBi7LR5eztDySbK5m+dj3pC7X6NCelMUpP3CYkhhjCYYbLqez2g
Mm7VPBO4sqdL4npbdC8I6A07V6SSDMK3vRltBiYtuJnHDrIEL9hkH2JTSktvIu0Y
/b51vo2v/GpYpaoGH0COIQFAokw9VYAevuoHCDEjdliVxFShvWvJm+rxTAg6JEUW
XuXmJ7LPOX6peJVNsR6n3BXiEGDmFS4qelxwXcoP4xI6J07XflZZWoj5pmdsbrj8
XgIjGfvJDh4sw5jy0BMeWl9qhP1NM+kpM4SYove6zV/WnPaAPbKgWPwxTZ0uXg+6
XQ3klGUHyQ3yc6J+AmBDnHM3/9tdIYtUsIPjMjlPjO/fuu+7y4vW++H0S7wXU2mE
UBR/uAKywT4dMbgKauCLxrirU7a+zPiABbvZnG9ItWaXsUjoTED1AaAR2shr3/ih
j8TifrDqmPFW4GyNvveaUTBGlQMj2CO6r/7FNem0ltcgMZh89uRWX2C9dGzrwHs0
WyUC/of9Ml1E2eW9uJdu2OdkN07YZ0r445TRPoycj8sqfCA86G4RAAZQowNc3KOh
gCGF8aKoWop/RdpgslGALnZViMBKF2WBgxU3hVsuqv/+O5g76Uj3+HR88Nv56ZNT
U0UN5CwLOGatHhubb5LuHzgNw25+0rwxu4sBSqdx2XLhZborwy//cVybVcnKEt8t
zOMedj2KLduzc9inIkc/eNFjBwndTBObGlAYJg/JIvMfka5dC1LTBgVTqYtAOfnH
bUPikEg2kMdtO+Sq28t9mhqodP5aajGom1aBXm+M3HNvqL83XrrnE57pzlA3pxo+
1FU2OQgXYq/D6FjhhRDzjy8xlIJwhhCm29vQL6uXdeEOj7WlVnjWOVsZlXn/bgIN
eNxXxy+fQkhF5QuZzrMtxz0zdGtEllscYqV1SjrP8nifDZCvT/YwmqVYR3zuaAat
g7Gn1adylV3dJZzuaE+rni1VHXflqD/03jlp4X4yh1/eZmG+4xSgdPPEIOQMkkaI
FuT+wVwZEDgC4RUWFSW/uqK+7qUz57NvAXulSDbvWZ1aliMYev81buKo3K1UxnWI
l9AhEuxuQPS9hMtHtCqeVLHhIHI1iq1I/tit85XoCOre9JtmoBBsVEOnkWDuGvQf
Cks2cZEHaNq6r1EwqcM5s1+ZuthAJKQ5HWz4nujPK8/QVuaYZ6KsEkI2c+bNebuz
HdGplUu1yXXpYCbssRCQzEemtyOt+B5J83LZV7Y45UlHhYC9Ss7QA3CFVTtFci9g
K1bAJhWGZUA81+wf3NA8nKmB8BUT1/v+51d5DUpKaWm/+e04TejbSVfM3g47ZICe
ybGUUG8dDuEWGo62pv2QOtiN3K5PvkiCBxf8zl1g8kbMzTzbQUIgggLgJMhmIz1a
VHaflUNdq2NV1KJ1W/TV7c+lD7Q2IUgnZYIVXlp1n841J3QYTN7Ms+X13/4QdwYh
tElOsINwFdZ3DMaTAPoSre411s5RgfjrueEP5A9Qb8xVwB1UQbdM0YAyB8CVfmBa
1PfpPg/9NA66lyj05Q/JBXkqVCxlqizJJKpAEgWB1C9RFdVCvdt3GhFX0NHbVE9y
HNtBqdkI9+ZxTyKet6ZmNIc82sBksDTsl3Lq8Q/1vIr4GxFxVWeaOiuf32v6Kwy7
hpbuPz1IBwqV+S64S9zviSahAfX4TEETQ9VLIUZLWyhPV/jZ/GBxQLWtW1O4VHF7
JQhBbATapANdBJjxrJ+7Xn7yoIHv7COkoSZyz/FSKLhBppmnSUkjHvn6QdSbETuV
rMfpu3iLX43i13PzDUPXHpJW+leWZLCdNVAXvpvAUn/ufOIErbv+K+trwbESzmuy
K5rLU9FoYQsvBlsq10oU13Xeu9xLfSLPApLbOBVjhCiz3kyxhpP8ufCP4A48nrVi
nvILWlCyI4lCTCc2HXRpOtM8ooyCSsXik/k1bTS0qVoZUerzXaQbhjuA9BMOA0Cw
9pWX6l7J3qsl6ovVEycZ+QY2m6xmV3FaLSk5JrOstdc3jp521tQM/8aYF5ejx8yW
z1P0zPF61dM2+1Zdx5ueY5+nDIo+Ri6sRXTu2fiQSBB55IPpbHIM/5+/bpclKaW8
5dusdlVLAJPPpEk+Qq0gGZMknYVY+hMWpJCk2oeuvNCdXaC4o0TITKAAB6HWTZaZ
0MM7+7F1Rdm1O+7URKfVZuUv+HSS218RaJW72IiEIV6dhuXHiyXgjkZEmiF0cl6F
HLXbgnfZaO3CBqp9R5B1ZaVryeveh6xoGev2rwYS4wuQtAIbcoKPTKAmxddGysKB
dnNErnOx/jFvpTbj17L89MWl9wJPoOpt/72FWtwxB6YhDXac3YXRikW91paU/eNw
XUu71y2CEUb8lL3QsBUWxsQRPttUbvZW8Yo6K6pLoYLLp4Z5+eupbPhquNBP1cgf
G9ssJWAZnMGBDO2QzKzAZU3QhM5tZq44MOX9h7rcUqMX4VRFf40ti9Tg4b8dn/BV
T6mVdmKYBM+6I1Q0K+H6sj+4MOIZQVSDfvt+ucZ9bXBWL6iJfLh8zSuc6KZaCqeu
VTys9+MI55CMt0QUq7edN8rvoNgjaiOaOHoR+pjCdieJedx8nxA5fBxYLO0aKEJS
GzLu0WafB8o9SAdEgLoxDClbUxV0SwrzYrjoXamzA6QyGXOEiAKIZSPvjJvmKRgm
BFv1XXNhQMUOWZhbIPTgNzh9spxAQa3ioVQtwr2NAO/a10vdrqY7Ej88h1DJA0+Q
LGzZmHGrz+Fx1m4XXS5jBidfyjPydZxPH84ga2t1JlsAHIBSQFFOUDQYj0sb+cp+
bvgoG1De/c2ijGb3+fPYNz9Wd0Erdgkd6nh77NQG/Sv+4iTAUBK9WTqLNBPci99b
pvAE169Lj5EBd4Zm/NGsogs2BW4kK9icF+zpSAaBa2/BYcVK2cN2BaXHKXuIIqD5
9k6vniLpleN636oS3s6mUTaO9zCiEiuS8DNmNbndcnac/rvx302ws5xJWk7wjo8s
lAGY8+8LMmDtg+1B+KVMBvvjJswOKKpBJbuOkSSFXYqwt55iHzPLmLAZbdOO8HmC
5XsUXwdbn1Pnvxb03sk9396DxJuwHerWmegx8BqkM2K/SEupj68UhWQ+i1sdq/GA
Y/p/k3/WO6NV45ekzpprY9ubl6BX9tkp3pyEsVV+1fliBC+yHC2dLZrfKJOYpL2F
66rw0I9ILbFScFZTWj52/CTI0P8F07bkaZ+/Wn/XvNMx8YoOh9xXTlEvDnaA+qMM
2EKgzPHV/FIjFhJn2WLjIrCcxlFyCfFbAuwD8a+GUHqUMYViohvo85Y4dUqLLUaD
FD492WXVcviJBw5pMnzYFPIYDDA6r2YHHGb8HjsJh8kn8lT2twneblv5ypuKqccn
BPyvJ/gttrLnVlPI3Pcc/+SD+u89x5kiJ2oEh42IE5K+dmvos5wGKi8aqv8C38Il
B8l2daxQoUJofH2InW9mXUHbVJ8vj8jDI9w2VvJMmFIzRnld8uN4siAxJ0/6my0I
3XBSiHunwnhtbEBQqaIe3V8yJ3kcMdF+zV7sNl74ciyrz/0zHGsPFK8ZEn7A8Tmn
Nk/os2TbRA29H4+7owFPIej09tcg0mju3lxkt3l8V3FVWJCUM2yzFsKr12Y+1b9g

//pragma protect end_data_block
//pragma protect digest_block
DoTMndGzG+hf3cY8wMpEA2iO8go=
//pragma protect end_digest_block
//pragma protect end_protected
